`include "../rf32x32.v"

module register_test;
  reg

  endmodule