module ifid(order_data, pc_out_data, plusFour_out_data)

inout [31:0] order_data;
inout [31:0] pc_out_data;
inout [31:0] plusFour_out_data;

endmodule